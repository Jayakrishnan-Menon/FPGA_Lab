module venmachm_tb;
  
  reg clk;
  reg rst;
  reg [1:0] coin;
  wire chocolate,chips,biscuit;

endmodule
